module Hot_Block_Ring_Counter();

endmodule
